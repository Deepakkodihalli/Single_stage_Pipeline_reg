module pipeline_reg (
    input  logic        clk,
    input  logic        rst,      
    input  logic [7:0]  in,
    input  logic        in_valid,
    output logic        in_ready,
    output logic [7:0]  out,
    output logic        out_valid,
    input  logic        out_ready
);

   
    assign in_ready = ~out_valid || out_ready;

    always_ff @(posedge clk) begin
        if (!rst) begin
            out_valid <= 1'b0;
            out       <= 8'b0;
        end
        else begin
           
            if (in_valid && in_ready) begin
                out       <= in;
                out_valid <= 1'b1;
            end
          
            else if (out_valid && out_ready) begin
                out_valid <= 1'b0;
            end
        end
    end

endmodule

